
module sysclkout (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
